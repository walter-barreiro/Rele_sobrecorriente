IDMT_SI_200_01_rom_inst : IDMT_SI_200_01_rom PORT MAP (
		address	 => address_sig,
		clock	 => clock_sig,
		q	 => q_sig
	);
