sqrt_wizard_inst : sqrt_wizard PORT MAP (
		radical	 => radical_sig,
		q	 => q_sig,
		remainder	 => remainder_sig
	);
