lpm_add_sub_wizard_inst : lpm_add_sub_wizard PORT MAP (
		add_sub	 => add_sub_sig,
		dataa	 => dataa_sig,
		datab	 => datab_sig,
		result	 => result_sig
	);
